
module TOP_eg ( 
	`ifdef USE_POWER_PINS
		inout vssa1,
		inout vdda1
	`endif
  );
  
endmodule

